//Test bench for halfsubtactor
`include "half_sub.v"

module testbench;
    reg a, b;
    wire inverse_a, diff, borrow;
    
endmodule