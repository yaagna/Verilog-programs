// Verilog program of 4 bit carry look ahead adder

module cla4(a, b, cin, cout, y);
    input [3:0] a, b;
    input cin;
    output cout;
    output [3:0] y;

endmodule