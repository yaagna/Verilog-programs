// Testbench for 4-bit ALU

`include "alu_4bit.v"

module testbench;

endmodule