module mux4_1(input [3:0] i, output y, input [1:0] s);

endmodule