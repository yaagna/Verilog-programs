//Test bench for sr latch
`include "sr_latch.v"

module testbench;


endmodule