module mux();
    input 
    output

endmodule
