// Verilog 1 to 2 Demultiplexer program

module demux1_2();
    

endmodule