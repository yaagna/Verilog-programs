`include "full_adder.v"

module testbench;
    reg a, b, cin;
    wire sum, cout;
    
endmodule