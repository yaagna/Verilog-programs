// 4 bit ALU using Verilog HDL

module alu();

endmodule