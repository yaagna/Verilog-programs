module jk_latch(j, k, clk, reset, q);

    input j, k, clk, reset;
    output reg q;

endmodule