// Test bench for 1 to 4 demultiplexer
`include "demux1_4.v"

module testbench;

endmodule