module mux();


endmodule
