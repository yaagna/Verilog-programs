// Test bench for 1 to 2 demultiplexer

module testbench;

endmodule

//iverilog -o demux1_2_testbench.vvp demux1_2_testbench.v
//vvp demux1_2_testbench.vvp
