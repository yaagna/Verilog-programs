//Testbench for JK latch
`include "jk_latch.v"

module testbench;
    

endmodule