// Verilog 1 to 4 Demultiplexer program using behavioural model

module demux1_4();

endmodule