module (i0, i1, s, y);
    input wire i0, i1, s;
    output y;

    

endmodule