//Testbench for JK latch
`include "jk_latch.v"

module testbench;
    reg j;
    reg k;
    reg clk;
    reg reset;
    output reg q;

    initial clk = 0;

endmodule